//Just a dummy module to try out the New trans_receiver module